LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

package Utiles is
	
	type genericArrayofVector16bit is array (natural range <>) of std_logic_vector(15 downto 0);


end Utiles;


-- Package Body Section
package body Utiles is

	
end Utiles;


